package spi_pkg;
  
    import uvm_pkg::*;
    import wb2spi_pkg::*;
    import wb2spi_parameters_pkg::*;
    `include "uvm_macros.svh"
    `include "timescale.v"
    `include "spi_macros.svh"
    `include "spi_defines.svh"
    `include "spi_transaction.svh"
    `include "spi_configuration.svh"
    `include "spi_driver.svh"
    `include "spi_monitor.svh"
    `include "spi_sequence_base.svh"
    `include "spi_agent.svh"

endpackage