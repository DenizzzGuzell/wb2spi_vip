package spi_pkg_hdl;
  `include "spi_macros.svh"
  `include "spi_defines.svh"
endpackage