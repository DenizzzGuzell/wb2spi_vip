package wb2spi_scoreboard_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"



    import wb_pkg::*;
    import spi_pkg::*;
    import wb2spi_env_cfg_pkg::*;
    `include "scoreboard_macros.svh"
    `include "wb2spi_scoreboard.svh"
endpackage