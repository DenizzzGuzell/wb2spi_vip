package wb2spi_parameters_pkg;

    parameter int SPI_SS_NB = 8;

    parameter string spi_BFM  = "spi_BFM";
    parameter string wb_BFM  = "wb_BFM";

    parameter string AGENT_CONFIGS = "AGENT_CONFIGS";
    parameter string CONFIGURATIONS = "CONFIGURATIONS";
    parameter string MONITORS = "MONITORS";
    parameter string SEQUENCERS = "SEQUENCERS";
    
endpackage