package wb2spi_env_cfg_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  //import spi_pkg::*;
  //import spi_pkg_hdl::*;
  import wb2spi_pkg::*;
  import wb_pkg::*;
  import wb_pkg_hdl::*;
  import spi_pkg::*;
  import spi_pkg_hdl::*;
  `include "timescale.v"
  `include "wb2spi_environment_configuration.svh"


endpackage