`include "timescale.v"
package wb2spi_pkg;

    `include "wb2spi_macros.svh"
    `include "timescale.v"

endpackage