package wb_pkg_hdl;
  
  `include "wb_macros.svh"

endpackage