package wb_pkg;
  
    import uvm_pkg::*;
    import wb2spi_pkg::*;
    import wb2spi_parameters_pkg::*;
    `include "uvm_macros.svh"
    `include "timescale.v"
    `include "wb_macros.svh"
    `include "wb_transaction.svh"
    `include "wb_configuration.svh"
    `include "wb_driver.svh"
    `include "wb_monitor.svh"
    `include "wb_sequence_base.svh"
    `include "wb2reg_adapter.svh"
    `include "wb_agent.svh"

endpackage