package wb2spi_tests_pkg;

   import uvm_pkg::*;
   import wb2spi_pkg::*;
   import wb2spi_parameters_pkg::*;
   import wb2spi_env_cfg_pkg::*;
   import wb2spi_env_pkg::*;
   import wb2spi_sequences_pkg::*;
   import wb_pkg::*;
   import wb_pkg_hdl::*;
   import spi_pkg::*;
   import spi_pkg_hdl::*;

   `include "uvm_macros.svh"
   `include "timescale.v"

   `include "wb2spi_test_base.svh"
   `include "wb2spi_example_test.svh"


endpackage